

module letterROMSV(
// input is the letter and the X and Y value on the specified region. If the letterrom array has 1 on that pixel then we enable write, o/w we don't
input [3:0] letter,	   // whether it is A,B,C...
input [7:0] x,					// xth pixel on screen 
input [6:0] y,					// yth pixel on screen
output pixel				// whether it is 1 or zero
);

// Each letter is represented by 8*16 pixels and since there are 16 letters we will have 8*(16 * 16) = 8 * 255 sized array

logic [0:7] letter_rom [0:255]=
'{
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00010000, // 2    *
		8'b00111000, // 3   ***
		8'b01101100, // 4  ** **
		8'b11000110, // 5 **   **
		8'b11000110, // 6 **   **
		8'b11111110, // 7 *******
		8'b11000110, // 8 **   **
		8'b11000110, // 9 **   **
		8'b11000110, // a **   **
		8'b11000110, // b **   **
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// B: 2
		8'b00000000, // 0
		8'b00000000, // 1
		8'b11111100, // 2 ******
		8'b01100110, // 3  **  **
		8'b01100110, // 4  **  **
		8'b01100110, // 5  **  **
		8'b01111100, // 6  *****
		8'b01100110, // 7  **  **
		8'b01100110, // 8  **  **
		8'b01100110, // 9  **  **
		8'b01100110, // a  **  **
		8'b11111100, // b ******
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// C: 3
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00111100, // 2   ****
		8'b01100110, // 3  **  **
		8'b11000010, // 4 **    *
		8'b11000000, // 5 **
		8'b11000000, // 6 **
		8'b11000000, // 7 **
		8'b11000000, // 8 **
		8'b11000010, // 9 **    *
		8'b01100110, // a  **  **
		8'b00111100, // b   ****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// D: 4
		8'b00000000, // 0
		8'b00000000, // 1
		8'b11111000, // 2 *****
		8'b01101100, // 3  ** **
		8'b01100110, // 4  **  **
		8'b01100110, // 5  **  **
		8'b01100110, // 6  **  **
		8'b01100110, // 7  **  **
		8'b01100110, // 8  **  **
		8'b01100110, // 9  **  **
		8'b01101100, // a  ** **
		8'b11111000, // b *****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// 5
		8'b00000000, // 0
		8'b00000000, // 1
		8'b11111110, // 2 *******
		8'b01100110, // 3  **  **
		8'b01100010, // 4  **   *
		8'b01101000, // 5  ** *
		8'b01111000, // 6  ****
		8'b01101000, // 7  ** *
		8'b01100000, // 8  **
		8'b01100010, // 9  **   *
		8'b01100110, // a  **  **
		8'b11111110, // b *******
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// 6
		8'b00000000, // 0
		8'b00000000, // 1
		8'b11111110, // 2 *******
		8'b01100110, // 3  **  **
		8'b01100010, // 4  **   *
		8'b01101000, // 5  ** *
		8'b01111000, // 6  ****
		8'b01101000, // 7  ** *
		8'b01100000, // 8  **
		8'b01100000, // 9  **
		8'b01100000, // a  **
		8'b11110000, // b ****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// 7
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00111100, // 2   ****
		8'b01100110, // 3  **  **
		8'b11000010, // 4 **    *
		8'b11000000, // 5 **
		8'b11000000, // 6 **
		8'b11011110, // 7 ** ****
		8'b11000110, // 8 **   **
		8'b11000110, // 9 **   **
		8'b01100110, // a  **  **
		8'b00111010, // b   *** *
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// H: 8
		8'b00000000, // 0
		8'b00000000, // 1
		8'b11000110, // 2 **   **
		8'b11000110, // 3 **   **
		8'b11000110, // 4 **   **
		8'b11000110, // 5 **   **
		8'b11111110, // 6 *******
		8'b11000110, // 7 **   **
		8'b11000110, // 8 **   **
		8'b11000110, // 9 **   **
		8'b11000110, // a **   **
		8'b11000110, // b **   **
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// I: 9
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00111100, // 2   ****
		8'b00011000, // 3    **
		8'b00011000, // 4    **
		8'b00011000, // 5    **
		8'b00011000, // 6    **
		8'b00011000, // 7    **
		8'b00011000, // 8    **
		8'b00011000, // 9    **
		8'b00011000, // a    **
		8'b00111100, // b   ****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// J: a
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00011110, // 2    ****
		8'b00001100, // 3     **
		8'b00001100, // 4     **
		8'b00001100, // 5     **
		8'b00001100, // 6     **
		8'b00001100, // 7     **
		8'b11001100, // 8 **  **
		8'b11001100, // 9 **  **
		8'b11001100, // a **  **
		8'b01111000, // b  ****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// K: b
		8'b00000000, // 0
		8'b00000000, // 1
		8'b11100110, // 2 ***  **
		8'b01100110, // 3  **  **
		8'b01100110, // 4  **  **
		8'b01101100, // 5  ** **
		8'b01111000, // 6  ****
		8'b01111000, // 7  ****
		8'b01101100, // 8  ** **
		8'b01100110, // 9  **  **
		8'b01100110, // a  **  **
		8'b11100110, // b ***  **
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// L: c
		8'b00000000, // 0
		8'b00000000, // 1
		8'b11110000, // 2 ****
		8'b01100000, // 3  **
		8'b01100000, // 4  **
		8'b01100000, // 5  **
		8'b01100000, // 6  **
		8'b01100000, // 7  **
		8'b01100000, // 8  **
		8'b01100010, // 9  **   *
		8'b01100110, // a  **  **
		8'b11111110, // b *******
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// M: d
		8'b00000000, // 0
		8'b00000000, // 1
		8'b11000110, // 2 **   **
		8'b11101110, // 3 *** ***
		8'b11111110, // 4 *******
		8'b11111110, // 5 *******
		8'b11010110, // 6 ** * **
		8'b11000110, // 7 **   **
		8'b11000110, // 8 **   **
		8'b11000110, // 9 **   **
		8'b11000110, // a **   **
		8'b11000110, // b **   **
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// N: e
		8'b00000000, // 0
		8'b00000000, // 1
		8'b11000110, // 2 **   **
		8'b11100110, // 3 ***  **
		8'b11110110, // 4 **** **
		8'b11111110, // 5 *******
		8'b11011110, // 6 ** ****
		8'b11001110, // 7 **  ***
		8'b11000110, // 8 **   **
		8'b11000110, // 9 **   **
		8'b11000110, // a **   **
		8'b11000110, // b **   **
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// O: f
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111100, // 2  *****
		8'b11000110, // 3 **   **
		8'b11000110, // 4 **   **
		8'b11000110, // 5 **   **
		8'b11000110, // 6 **   **
		8'b11000110, // 7 **   **
		8'b11000110, // 8 **   **
		8'b11000110, // 9 **   **
		8'b11000110, // a **   **
		8'b01111100, // b  *****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// P: code x50
		8'b00000000, // 0
		8'b00000000, // 1
		8'b11111100, // 2 ******
		8'b01100110, // 3  **  **
		8'b01100110, // 4  **  **
		8'b01100110, // 5  **  **
		8'b01111100, // 6  *****
		8'b01100000, // 7  **
		8'b01100000, // 8  **
		8'b01100000, // 9  **
		8'b01100000, // a  **
		8'b11110000, // b ****
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000 // f
};

assign pixel = letter_rom[16*letter +y][x];

endmodule